PASSED::tran L
VS 1 0 1 CONSTANT(1 0 1)
R1 1 2 1
L1 2 0 1N
.TRAN 0.1NS 20NS
.PLOT TRAN V(2)
.END