testing stamp utility 1: pure negative elements

R1 1 0 5
R2 1 2 6
VIN 2 0 DC 2

.DC VIN 0 5 0.1
.END
