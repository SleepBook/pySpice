Single Ressitor and Source

R1 1 0 20K
R2 1 2 2M
VIN 2 0 DC 6

.END
