testing stamping utility 2: xcxs

VIN 1 0 2
*I0 1 0 2
R1 1 2 10
E1 2 0 1 0 5

.DC VIN 0 5 0.1
.END