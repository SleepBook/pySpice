test stamping utility: ac and tran

VIN 1 0 DC 1 AC 1 SIN(0 10 300X)
C1 1 2 2
L1 2 0 3

.AC DEC 3 1 10K
.TRAN 1NS 100NS
.END